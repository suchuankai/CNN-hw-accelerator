`include "PE.v"
`include "PE_array.v"
`include "RfTemp.v"
`include "Adder.v"
`include "Adder2.v"
`include "psumBuf.v"
`include "convBuf.v"
`include "controller.v"
`include "FIFO.v"
`include "rowRf.v"
`include "rowSelect.v"
`include "FIFO_out.v"
`include "FIFO_w.v"
`include "demux1_3.v"
`include "biasBuf.v"
`include "weightBuf.v"
